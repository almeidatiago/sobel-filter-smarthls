-- ----------------------------------------------------------------------------
-- Smart High-Level Synthesis Tool Version 2021.1.2
-- Copyright (c) 2015-2021 Microchip Technology Inc. All Rights Reserved.
-- For support, please contact: smarthls@microchip.com
-- Date: Tue Nov 16 16:39:41 2021
-- ----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

-- SmartHLS generic types
package legup_types_pkg is
type slv_array_t is array (natural range <> ) of std_logic_vector;

end package legup_types_pkg;

package body legup_types_pkg is
end package body legup_types_pkg;
